* File: OAI.pex.sp
* Created: Wed Oct 26 07:31:45 2022
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "OAI.pex.sp.pex"
.subckt OAI  OUT GND! VDD! D C A B
* 
* B	B
* A	A
* C	C
* D	D
* VDD!	VDD!
* GND!	GND!
* OUT	OUT
XD0_noxref N_GND!_D0_noxref_pos N_VDD!_D0_noxref_neg DIODENWX  AREA=9.69563e-12
+ PERIM=1.2474e-05
XMMN2 N_OUT_MMN2_d N_D_MMN2_g N_NET17_MMN2_s N_GND!_D0_noxref_pos NFET L=7e-08
+ W=1e-06 AD=4.69e-13 AS=2.6e-13 PD=1.938e-06 PS=2.52e-06 NRD=0.325 NRS=0.1 M=1
+ NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=2.6e-07 SB=1.98e-06 SD=0 PANW1=0
+ PANW2=0 PANW3=7e-16 PANW4=3.5e-15 PANW5=3.5e-15 PANW6=7e-15 PANW7=1.4e-14
+ PANW8=1.4e-14 PANW9=2.73e-14 PANW10=0
XMMN3 N_OUT_MMN2_d N_C_MMN3_g N_NET17_MMN3_s N_GND!_D0_noxref_pos NFET L=7e-08
+ W=1e-06 AD=4.69e-13 AS=2.205e-13 PD=1.938e-06 PS=1.441e-06 NRD=0.613 NRS=0.102
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.268e-06 SB=9.72e-07 SD=0
+ PANW1=0 PANW2=0 PANW3=7e-16 PANW4=3.5e-15 PANW5=3.5e-15 PANW6=7e-15
+ PANW7=1.4e-14 PANW8=1.4e-14 PANW9=2.73e-14 PANW10=0
XMMN0 N_NET17_MMN3_s N_A_MMN0_g N_GND!_MMN0_s N_GND!_D0_noxref_pos NFET L=7e-08
+ W=1e-06 AD=2.205e-13 AS=1.045e-13 PD=1.441e-06 PS=1.209e-06 NRD=0.339
+ NRS=0.107 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.779e-06
+ SB=4.61e-07 SD=0 PANW1=0 PANW2=0 PANW3=7e-16 PANW4=3.5e-15 PANW5=3.5e-15
+ PANW6=7e-15 PANW7=1.4e-14 PANW8=1.4e-14 PANW9=2.73e-14 PANW10=0
XMMN1 N_NET17_MMN1_d N_B_MMN1_g N_GND!_MMN0_s N_GND!_D0_noxref_pos NFET L=7e-08
+ W=1e-06 AD=1.82e-13 AS=1.045e-13 PD=2.364e-06 PS=1.209e-06 NRD=0.104 NRS=0.102
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=2.058e-06 SB=1.82e-07 SD=0
+ PANW1=0 PANW2=0 PANW3=7e-16 PANW4=3.5e-15 PANW5=3.5e-15 PANW6=7e-15
+ PANW7=1.4e-14 PANW8=1.4e-14 PANW9=2.73e-14 PANW10=0
XMMP3 NET15 N_D_MMP3_g N_VDD!_MMP3_s N_VDD!_D0_noxref_neg PFET L=7e-08 W=2e-06
+ AD=9.38e-13 AS=5.14e-13 PD=2.938e-06 PS=4.514e-06 NRD=0.2345 NRS=0.05 M=1 NF=1
+ CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.57e-07 SB=1.972e-06 SD=0 PANW1=0
+ PANW2=2.73e-15 PANW3=3.5e-15 PANW4=3.5e-15 PANW5=3.5e-15 PANW6=7e-15
+ PANW7=1.1148e-13 PANW8=8.2e-14 PANW9=5.6e-14 PANW10=8.4e-14
XMMP0 N_OUT_MMP0_d N_C_MMP0_g NET15 N_VDD!_D0_noxref_neg PFET L=7e-08 W=2e-06
+ AD=4.41e-13 AS=9.38e-13 PD=2.441e-06 PS=2.938e-06 NRD=0.051 NRS=0.2345 M=1
+ NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.265e-06 SB=9.64e-07 SD=0
+ PANW1=0 PANW2=2.73e-15 PANW3=3.5e-15 PANW4=3.5e-15 PANW5=3.5e-15 PANW6=7e-15
+ PANW7=2.548e-14 PANW8=2.8e-14 PANW9=5.6e-14 PANW10=3.64e-13
XMMP1 N_OUT_MMP0_d N_A_MMP1_g NET20 N_VDD!_D0_noxref_neg PFET L=7e-08 W=2e-06
+ AD=4.41e-13 AS=2.09e-13 PD=2.441e-06 PS=2.209e-06 NRD=0.1695 NRS=0.05225 M=1
+ NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.776e-06 SB=4.53e-07 SD=0
+ PANW1=0 PANW2=2.73e-15 PANW3=3.5e-15 PANW4=3.5e-15 PANW5=3.5e-15 PANW6=7e-15
+ PANW7=2.548e-14 PANW8=1.4e-13 PANW9=8.4e-14 PANW10=8.4e-14
XMMP2 NET20 N_B_MMP2_g N_VDD!_MMP2_s N_VDD!_D0_noxref_neg PFET L=7e-08 W=2e-06
+ AD=2.09e-13 AS=3.48e-13 PD=2.209e-06 PS=4.348e-06 NRD=0.05225 NRS=0.054 M=1
+ NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.055e-06 SB=1.74e-07 SD=0
+ PANW1=0 PANW2=2.73e-15 PANW3=3.5e-15 PANW4=3.5e-15 PANW5=3.5e-15 PANW6=7e-15
+ PANW7=1.6548e-13 PANW8=2.8e-14 PANW9=5.6e-14 PANW10=8.4e-14
c_243 NET15 0 2.66343e-19
*
.include "OAI.pex.sp.OAI.pxi"
*
.ends
*
*
