* File: AOAI211.pex.sp
* Created: Wed Oct 26 07:49:51 2022
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "AOAI211.pex.sp.pex"
.subckt AOAI211  GND! OUT VDD! D C A B
* 
* B	B
* A	A
* C	C
* D	D
* VDD!	VDD!
* OUT	OUT
* GND!	GND!
XD0_noxref N_GND!_D0_noxref_pos N_VDD!_D0_noxref_neg DIODENWX  AREA=9.69563e-12
+ PERIM=1.2474e-05
XMMN3 N_noxref_20_MMN3_d N_D_MMN3_g N_GND!_MMN3_s N_GND!_D0_noxref_pos NFET
+ L=7e-08 W=1e-06 AD=4.69e-13 AS=2.65e-13 PD=1.938e-06 PS=2.53e-06 NRD=0.62
+ NRS=0.1 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=2.65e-07 SB=1.971e-06
+ SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=9.1e-16 PANW5=3.5e-15 PANW6=7e-15
+ PANW7=1.4e-14 PANW8=1.4e-14 PANW9=2.8e-14 PANW10=2.59e-15
XMMN2 N_OUT_MMN2_d N_C_MMN2_g N_noxref_20_MMN3_d N_GND!_D0_noxref_pos NFET
+ L=7e-08 W=1e-06 AD=2.205e-13 AS=4.69e-13 PD=1.441e-06 PS=1.938e-06 NRD=0.102
+ NRS=0.318 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.273e-06
+ SB=9.63e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=9.1e-16 PANW5=3.5e-15
+ PANW6=7e-15 PANW7=1.4e-14 PANW8=1.4e-14 PANW9=2.8e-14 PANW10=2.59e-15
XMMN0 N_OUT_MMN2_d N_A_MMN0_g noxref_22 N_GND!_D0_noxref_pos NFET L=7e-08
+ W=1e-06 AD=2.205e-13 AS=1.045e-13 PD=1.441e-06 PS=1.209e-06 NRD=0.339
+ NRS=0.1045 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.784e-06
+ SB=4.52e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=9.1e-16 PANW5=3.5e-15
+ PANW6=7e-15 PANW7=1.4e-14 PANW8=1.4e-14 PANW9=2.8e-14 PANW10=2.59e-15
XMMN1 noxref_22 N_B_MMN1_g N_noxref_20_MMN1_s N_GND!_D0_noxref_pos NFET L=7e-08
+ W=1e-06 AD=1.045e-13 AS=1.73e-13 PD=1.209e-06 PS=2.346e-06 NRD=0.1045
+ NRS=0.104 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=2.063e-06
+ SB=1.73e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=9.1e-16 PANW5=3.5e-15
+ PANW6=7e-15 PANW7=1.4e-14 PANW8=1.4e-14 PANW9=2.8e-14 PANW10=2.59e-15
XMMP3 N_OUT_MMP3_d N_D_MMP3_g N_VDD!_MMP3_s N_VDD!_D0_noxref_neg PFET L=7e-08
+ W=2e-06 AD=9.38e-13 AS=5.14e-13 PD=2.938e-06 PS=4.514e-06 NRD=0.31 NRS=0.05
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.57e-07 SB=1.972e-06 SD=0
+ PANW1=0 PANW2=2.17e-15 PANW3=3.5e-15 PANW4=3.5e-15 PANW5=3.5e-15 PANW6=7e-15
+ PANW7=1.1204e-13 PANW8=8.2e-14 PANW9=5.6e-14 PANW10=8.4e-14
XMMP2 N_OUT_MMP3_d N_C_MMP2_g N_NET19_MMP2_s N_VDD!_D0_noxref_neg PFET L=7e-08
+ W=2e-06 AD=9.38e-13 AS=4.41e-13 PD=2.938e-06 PS=2.441e-06 NRD=0.159 NRS=0.051
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.265e-06 SB=9.64e-07 SD=0
+ PANW1=0 PANW2=2.17e-15 PANW3=3.5e-15 PANW4=3.5e-15 PANW5=3.5e-15 PANW6=7e-15
+ PANW7=2.604e-14 PANW8=2.8e-14 PANW9=5.6e-14 PANW10=3.64e-13
XMMP0 N_NET19_MMP2_s N_A_MMP0_g N_VDD!_MMP0_s N_VDD!_D0_noxref_neg PFET L=7e-08
+ W=2e-06 AD=4.41e-13 AS=2.09e-13 PD=2.441e-06 PS=2.209e-06 NRD=0.1695 NRS=0.052
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.776e-06 SB=4.53e-07 SD=0
+ PANW1=0 PANW2=2.17e-15 PANW3=3.5e-15 PANW4=3.5e-15 PANW5=3.5e-15 PANW6=7e-15
+ PANW7=2.604e-14 PANW8=1.4e-13 PANW9=8.4e-14 PANW10=8.4e-14
XMMP1 N_NET19_MMP1_d N_B_MMP1_g N_VDD!_MMP0_s N_VDD!_D0_noxref_neg PFET L=7e-08
+ W=2e-06 AD=3.48e-13 AS=2.09e-13 PD=4.348e-06 PS=2.209e-06 NRD=0.054 NRS=0.0525
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.055e-06 SB=1.74e-07 SD=0
+ PANW1=0 PANW2=2.17e-15 PANW3=3.5e-15 PANW4=3.5e-15 PANW5=3.5e-15 PANW6=7e-15
+ PANW7=1.6604e-13 PANW8=2.8e-14 PANW9=5.6e-14 PANW10=8.4e-14
*
.include "AOAI211.pex.sp.AOAI211.pxi"
*
.ends
*
*
