* File: INV.pex.SP
* Created: Wed Oct 26 07:13:01 2022
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "INV.pex.SP.pex"
.subckt INV  GND! OUT VDD! IN
* 
* IN	IN
* VDD!	VDD!
* OUT	OUT
* GND!	GND!
XD0_noxref N_GND!_D0_noxref_pos N_VDD!_D0_noxref_neg DIODENWX  AREA=5.09242e-12
+ PERIM=9.35e-06
XMMN4 N_OUT_MMN4_d N_IN_MMN4_g N_GND!_MMN4_s N_GND!_D0_noxref_pos NFET L=7e-08
+ W=1e-06 AD=2.7e-13 AS=2.65e-13 PD=2.54e-06 PS=2.53e-06 NRD=0.102 NRS=0.1 M=1
+ NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=2.65e-07 SB=2.7e-07 SD=0 PANW1=0
+ PANW2=0 PANW3=0 PANW4=9.1e-16 PANW5=3.5e-15 PANW6=7e-15 PANW7=1.4e-14
+ PANW8=1.4e-14 PANW9=2.8e-14 PANW10=2.59e-15
XMMP4 N_OUT_MMP4_d N_IN_MMP4_g N_VDD!_MMP4_s N_VDD!_D0_noxref_neg PFET L=7e-08
+ W=2e-06 AD=5.34e-13 AS=5.14e-13 PD=4.534e-06 PS=4.514e-06 NRD=0.051 NRS=0.05
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.57e-07 SB=2.67e-07 SD=0
+ PANW1=0 PANW2=2.17e-15 PANW3=3.5e-15 PANW4=3.5e-15 PANW5=3.5e-15 PANW6=7e-15
+ PANW7=1.1204e-13 PANW8=2.22e-13 PANW9=5.6e-14 PANW10=8.4e-14
*
.include "INV.pex.SP.INV.pxi"
*
.ends
*
*
